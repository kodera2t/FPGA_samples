module and_comb(A, B, Y);
input A, B;
output Y;
assign Y=A&B;
endmodule